module segBdec
(
	input [3:0] D,
	output segB
);

  //////////////////////////////////////////
  // Declare any needed internal signals //
  ////////////////////////////////////////
  reg [0:15] truth_table = 16'b0000_0110_00xx_xxxx;
  
  //////////////////////////////////////////////////////
  // Write STRUCTURAL verilog to implement segment B //
  ////////////////////////////////////////////////////
  assign segB = truth_table[D];

  
endmodule
